p1_1.cir
.TITLE Problem 1 - common mode gain

V1  2   0   SIN(0 5MV 1KHZ)
V2  4   0   SIN(0 5MV 1KHZ)
M1  3   2   1   1   NFET
M2  5   4   1   1   NFET
.MODEL NFET NMOS (KP=400U VTO=1)
RSS 1   7   62K
RD1 3   6   62K
RD2 5   6   62K
VDD 6   0   DC  15V
VSS 7   0   DC  -15V

.TRAN   10NS    1MS
.MEASURE TRAN vpp1 PP V(2)
.MEASURE TRAN vpp2 PP V(3)
.MEASURE TRAN common_gain param='vpp2/vpp1'

.PROBE
.END

p3.cir
.TITLE Problem 3

Vi  1   0   SIN(0 10V 1000HZ)
C1  0   1   0.1U
R1  0   1   1073
R2  1   2   1073
C2  2   3   0.22U
R4  3   4   10K
R3  4   0   6875
X1  4   1   3   OPAMP1

.SUBCKT OPAMP1  1   2   6
RIN     1   2   10MEG
EGAIN   3   0   1   2   100K
RP1     3   4   1K
CP1     4   0   1.5915UF
EBUFFER 5   0   4   0   1
ROUT    5   6   10
.ENDS

.TRAN   10NS    2MS
.MEASURE TRAN vo PP par('V(3)/2')
.PRINT TRAN V(3)
.PROBE
.END


Extra 1
.TITLE Simulation of JFET
V1 1 0 SIN(0 10 1KHZ)
R1 1 2 100
RG1 2 3 1.9M
RG2 2 0 0.6M
J1 4 2 0 JM1
.MODEL JM1 NJF IS=8N
VDD 3 0 DC 20V
RD 4 3 5K
C2 4 5 1
RL 5 0 10K

.TRAN   100NS    2MS
.PRINT TRAN V(5)

.MEASURE TRAN vpp PP V(5)

.PROBE
.END

Circuit_1

.TITLE Simulation of problem 1

V1		2		0		SIN(0 0.25 1KHZ)
V2		4		0		SIN(0 -0.25 1KHZ)
M1		3		2		1		0		NFET
M2		5		4		1		0		NFET

.MODEL NFET NMOS

RSS		1		7		75K
RD1		3		6		75K
RD2		5		6		75K

VDD		6		0		DC		15V
VSS		7		0		DC		-15V

.TRAN   100NS    2MS

*.SAVE TRAN VM(2) VM(4)
.MEASURE TRAN vpp1 PP V(2)
.MEASURE TRAN vpp2 PP par('V(3)-V(5)')
.MEASURE TRAN diff_gain param='vpp2/vpp1'



.PROBE
.END
